dean@freud.762:1412005523