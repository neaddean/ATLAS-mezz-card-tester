dean@freud.444:1398263295