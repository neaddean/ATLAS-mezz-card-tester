library IEEE;
use IEEE.STD_LOGIC_1164.all;

package common is

  type multi_array is array (integer range 3 downto 0) of std_logic_vector (7 downto 0);

end common;
